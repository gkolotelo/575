--------------------------------------------------
-- Laboratorio de Circuitos Logicos - Turma A   --
--------------------------------------------------
-- 135964 Guilherme Kairalla Kolotelo           --
-- 137943 Alexandre Seidy Ioshisaqui            --
--------------------------------------------------
-- Laboratorio 5: Timers e Relogios de          --
--                  Tempo Real                  --
--------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_signed.all;
use ieee.numeric_std;

entity counter_k is
    generic (
        -- Change 'n' for larger (or shorter) maximum values for 'k'
        n : natural := 8
    );
    port (
        -- Standard maximum value = (255)decimal = (11111111)binary
        k       : in natural;
        clock   : in STD_LOGIC;
        reset_n : in STD_LOGIC;
        Q       : out STD_LOGIC_VECTOR(n-1 downto 0)
    );
end entity;
architecture rtl of counter_k is
    signal k_bin: std_logic_vector(n-1 downto 0);
begin
    -- Converts natural input 'k' into binary vector of 'n' bits
    k_bin <= conv_std_logic_vector(k, n);
    PROCESS(clock, reset_n)
        variable value : std_logic_vector(n-1 downto 0);
        begin
            if (reset_n = '0') then
                -- initialize all bits with zeros
                value := (OTHERS => '0');
            elsif (rising_edge(clock)) then
                -- Counts until 'k', then resets.
                if (numeric_std.to_integer(numeric_std.unsigned(value)) < numeric_std.to_integer(numeric_std.unsigned(k_bin))) then
                    value := value + '1';
                else
                    value := (OTHERS => '0');
                end if;
            end if;
        Q <= value;
    end process;
end rtl;