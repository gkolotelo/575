LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY Exp1c IS
	PORT ( SW : IN STD_LOGIC_VECTOR(17 DOWNTO 0); 
			LEDR : OUT STD_LOGIC_VECTOR(17 DOWNTO 0)); -- red LEDs 
END Exp1c;





architecture mux_5to1 OF Exp1c IS
	component mux2to1
	port (a, b, s: in std_logic;
		m: out std_logic);
	end component mux2to1;
	
	signal u, v, w, x, y, o1, o2, o3, m: std_logic;
	signal s: std_LOGIC_VECTOR(2 downto 0);

begin
	u <= SW(0);
	v <= SW(1);
	w <= SW(2);
	x <= SW(3);
	y <= SW(4);
	
	LEDR(17 downto 15) <= SW(17 downto 15);
	LEDR(4 downto 0) <= SW(4 dowNTO 0);
	
	mux1: mux2to1 port map (u, v, SW(17), o1);
	mux2: mux2to1 port map (w, x, SW(17), o2);
	mux3: mux2to1 port map (o1, o2, SW(16), o3);
	mux4: mux2to1 port map (o3, y, SW(15), LEDR(9));

	
	
end mux_5to1;